#Comentario
Int idade ;
Int altura -> 23 ;
String nome ;
String rg -> "CNH" ;

 If 12 == 12
     Read idade ;
 end 

Repeat 5
    Write "oi" ;
end 
