#Comentario
Int idade ;
String Nome -> "Gabriel Oliveira";
If ( 1 == 1 )
    Repeat 4
        Write "Meu nome";
    end
    Read nome ;
end ;