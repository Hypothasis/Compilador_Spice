Int idade -> 123 ;
String nome -> "Gabriel" ;
String RG ;