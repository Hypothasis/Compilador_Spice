#Comentario
Int idade ;
String Nome -> "Gabriel Oliveira" ;

If 12 == 12
    Read idade ;
end ;

Repeat 4
    Write "Meu nome" ;
end ;


