->
!=
==
||
&&
;
+
-
*
/
#Comentario
,
(
)