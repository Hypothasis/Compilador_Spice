Int idade ;
String nome ;