Int b;
Int a;