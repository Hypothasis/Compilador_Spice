;
Int abc ;
String bcd ;