#Declarando Inteiro, Inicializando e Atribuindo
Int idade ;
Int altura -> 1 ;
idade -> 21 ;

#Declarando String, Inicializando e Atribuindo
String nome ;
String RG -> "CNH" ;
nome -> "Gabriel" ;

#If
If 12 == 12
     Read idade ;
end 

#Repeat
Repeat 5
    Write "oi" ;
end 
